module not_gate (o1,i1);
input i1;
output o1;
not (o1,i1);
endmodule 