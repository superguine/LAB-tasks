module or_gate (o1,i1,i2);
input i1,i2;
output o1;
or (o1,i1,i2);
endmodule 